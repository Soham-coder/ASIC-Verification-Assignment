import uvm_pkg::*;
`include "uvm_macros.svh"
//`include "ASIC_config_obj.svh"
`include "definition_pkg.sv"
import definitions :: *;
`include "packet.sv"
`include "driver.sv"
`include "monitor.sv"
`include "sequencer.sv"
`include "packet_seqs.sv"
`include "agent.sv"
`include "env.sv"
`include "test_lib.sv"